module tables
(
	input rst_n,
	input [5:0] index,
	output [15:0] qe_out,
	output [5:0] nmps_out,
	output [5:0] nlps_out,
	output switch_out
);


reg [15:0] qe[0:46];
reg [5:0] nmps[0:46];
reg [5:0] nlps[0:46];
reg switch[0:46];

assign qe_out=qe[index];
assign nmps_out=nmps[index];
assign nlps_out=nlps[index];
assign switch_out=switch[index];
//初始化查找表
always @(negedge rst_n)
	if(!rst_n)begin
		qe[0]<=16'd22017;
		qe[1]<=16'd13313;
		qe[2]<=16'd6145;
		qe[3]<=16'd2753;
		qe[4]<=16'd1313;
		qe[5]<=16'd545;
		qe[6]<=16'd22017;
		qe[7]<=16'd21505;
		qe[8]<=16'd18433;
		qe[9]<=16'd14337;
		qe[10]<=16'd12289;
		qe[11]<=16'd9217;
		qe[12]<=16'd7169;
		qe[13]<=16'd5633;
		qe[14]<=16'd22017;
		qe[15]<=16'd21505;
		qe[16]<=16'd20737;
		qe[17]<=16'd18433;
		qe[18]<=16'd14337;
		qe[19]<=16'd13313;
		qe[20]<=16'd12289;
		qe[21]<=16'd10241;
		qe[22]<=16'd9217;
		qe[23]<=16'd8705;
		qe[24]<=16'd7169;
		qe[25]<=16'd6145;
		qe[26]<=16'd5633;
		qe[27]<=16'd5121;
		qe[28]<=16'd4609;
		qe[29]<=16'd4353;
		qe[30]<=16'd2753;
		qe[31]<=16'd2497;
		qe[32]<=16'd2209;
		qe[33]<=16'd1313;
		qe[34]<=16'd1089;
		qe[35]<=16'd673;
		qe[36]<=16'd545;
		qe[37]<=16'd321;
		qe[38]<=16'd273;
		qe[39]<=16'd133;
		qe[40]<=16'd73;
		qe[41]<=16'd37;
		qe[42]<=16'd21;
		qe[43]<=16'd9;
		qe[44]<=16'd5;
		qe[45]<=16'd1;
		qe[46]<=16'd22017;
		switch[0]<=1'd1;
		switch[1]<=1'd0;
		switch[2]<=1'd0;
		switch[3]<=1'd0;
		switch[4]<=1'd0;
		switch[5]<=1'd0;
		switch[6]<=1'd1;
		switch[7]<=1'd0;
		switch[8]<=1'd0;
		switch[9]<=1'd0;
		switch[10]<=1'd0;
		switch[11]<=1'd0;
		switch[12]<=1'd0;
		switch[13]<=1'd0;
		switch[14]<=1'd1;
		switch[15]<=1'd0;
		switch[16]<=1'd0;
		switch[17]<=1'd0;
		switch[18]<=1'd0;
		switch[19]<=1'd0;
		switch[20]<=1'd0;
		switch[21]<=1'd0;
		switch[22]<=1'd0;
		switch[23]<=1'd0;
		switch[24]<=1'd0;
		switch[25]<=1'd0;
		switch[26]<=1'd0;
		switch[27]<=1'd0;
		switch[28]<=1'd0;
		switch[29]<=1'd0;
		switch[30]<=1'd0;
		switch[31]<=1'd0;
		switch[32]<=1'd0;
		switch[33]<=1'd0;
		switch[34]<=1'd0;
		switch[35]<=1'd0;
		switch[36]<=1'd0;
		switch[37]<=1'd0;
		switch[38]<=1'd0;
		switch[39]<=1'd0;
		switch[40]<=1'd0;
		switch[41]<=1'd0;
		switch[42]<=1'd0;
		switch[43]<=1'd0;
		switch[44]<=1'd0;
		switch[45]<=1'd0;
		switch[46]<=1'd0;
		nmps[0]<=6'd1;
		nmps[1]<=6'd2;
		nmps[2]<=6'd3;
		nmps[3]<=6'd4;
		nmps[4]<=6'd5;
		nmps[5]<=6'd38;
		nmps[6]<=6'd7;
		nmps[7]<=6'd8;
		nmps[8]<=6'd9;
		nmps[9]<=6'd10;
		nmps[10]<=6'd11;
		nmps[11]<=6'd12;
		nmps[12]<=6'd13;
		nmps[13]<=6'd29;
		nmps[14]<=6'd15;
		nmps[15]<=6'd16;
		nmps[16]<=6'd17;
		nmps[17]<=6'd18;
		nmps[18]<=6'd19;
		nmps[19]<=6'd20;
		nmps[20]<=6'd21;
		nmps[21]<=6'd22;
		nmps[22]<=6'd23;
		nmps[23]<=6'd24;
		nmps[24]<=6'd25;
		nmps[25]<=6'd26;
		nmps[26]<=6'd27;
		nmps[27]<=6'd28;
		nmps[28]<=6'd29;
		nmps[29]<=6'd30;
		nmps[30]<=6'd31;
		nmps[31]<=6'd32;
		nmps[32]<=6'd33;
		nmps[33]<=6'd34;
		nmps[34]<=6'd35;
		nmps[35]<=6'd36;
		nmps[36]<=6'd37;
		nmps[37]<=6'd38;
		nmps[38]<=6'd39;
		nmps[39]<=6'd40;
		nmps[40]<=6'd41;
		nmps[41]<=6'd42;
		nmps[42]<=6'd43;
		nmps[43]<=6'd44;
		nmps[44]<=6'd45;
		nmps[45]<=6'd45;
		nmps[46]<=6'd46;
		nlps[0]<=6'd1;
		nlps[1]<=6'd6;
		nlps[2]<=6'd9;
		nlps[3]<=6'd12;
		nlps[4]<=6'd29;
		nlps[5]<=6'd33;
		nlps[6]<=6'd6;
		nlps[7]<=6'd14;
		nlps[8]<=6'd14;
		nlps[9]<=6'd14;
		nlps[10]<=6'd17;
		nlps[11]<=6'd18;
		nlps[12]<=6'd20;
		nlps[13]<=6'd21;
		nlps[14]<=6'd14;
		nlps[15]<=6'd14;
		nlps[16]<=6'd15;
		nlps[17]<=6'd16;
		nlps[18]<=6'd17;
		nlps[19]<=6'd18;
		nlps[20]<=6'd19;
		nlps[21]<=6'd19;
		nlps[22]<=6'd20;
		nlps[23]<=6'd21;
		nlps[24]<=6'd22;
		nlps[25]<=6'd23;
		nlps[26]<=6'd24;
		nlps[27]<=6'd25;
		nlps[28]<=6'd26;
		nlps[29]<=6'd27;
		nlps[30]<=6'd28;
		nlps[31]<=6'd29;
		nlps[32]<=6'd30;
		nlps[33]<=6'd31;
		nlps[34]<=6'd32;
		nlps[35]<=6'd33;
		nlps[36]<=6'd34;
		nlps[37]<=6'd35;
		nlps[38]<=6'd36;
		nlps[39]<=6'd37;
		nlps[40]<=6'd38;
		nlps[41]<=6'd39;
		nlps[42]<=6'd40;
		nlps[43]<=6'd41;
		nlps[44]<=6'd42;
		nlps[45]<=6'd43;
		nlps[46]<=6'd46;
	end

		

endmodule 