`timescale 1ns/1ns
module testbench3();



reg [7:0] data=8'd261;

wire data0=data[0];
wire data1=data[1];
wire data2=data[2];
wire data3=data[3];
wire data4=data[4];
wire data5=data[5];
wire data6=data[6];
wire data7=data[7];


endmodule 