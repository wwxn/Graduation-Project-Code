library verilog;
use verilog.vl_types.all;
entity code_queue_tb is
end code_queue_tb;
